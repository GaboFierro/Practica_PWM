module cycle_counter();